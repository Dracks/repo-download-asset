module github

pub struct Project {
	owner string [required]
	project string [required]
}